module clk_tree(
input wire in,
output out0,
output out1);

assign out0 = in;
assign out1 = in;


endmodule
