module clk_tree(
input wire in,
output out0,
output out1,
output out2,
output out3);

assign out0 = in;
assign out1 = in;
assign out2 = in;
assign out3 = in;

endmodule
